module crossbar();


endmodule