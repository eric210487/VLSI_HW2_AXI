module arbitration(

);
endmodule
module decoder(

);
endmodule