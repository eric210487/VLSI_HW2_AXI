module sram_wrapper(

);
endmodule